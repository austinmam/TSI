*MCP600X Comparator Test
.include C:\Users\nessa\Desktop\TSI\SPICE_subcircuits\MCP6001.sub
*.SUBCKT MCP6001 1 2 3 4 5
*                | | | | |
*                | | | | Output
*                | | | Negative Supply
*                | | Positive Supply
*                | Inverting Input
*                Non-inverting Input
*

Vcc Vcc 0 DC 5

Vpos Vpos 0 DC 5
Vneg Vneg 0 DC 2.5

X1 Vpos Vneg Vcc 0 Vout MCP6001

.DC Vpos 0 5.0 0.01

.probe
.end