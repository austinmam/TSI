* C:\Users\nessa\Desktop\TSI\ThrottlePlausibility\ThrottlePlausibility.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 2/16/2017 2:59:51 PM

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
R5  +10V Net-_R5-Pad2_ 1000		
R7  Net-_R6-Pad2_ RTN_+5V_ 1000		
R6  Net-_R5-Pad2_ Net-_R6-Pad2_ 8000		
R8  +5V Net-_R8-Pad2_ 1000		
R10  Net-_R10-Pad1_ GND 1000		
R9  Net-_R8-Pad2_ Net-_R10-Pad1_ 8000		
U1  Net-_R4-Pad1_ Net-_R2-Pad1_ Net-_R1-Pad1_ +5V Net-_R11-Pad2_ Net-_R4-Pad1_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_R12-Pad2_ Net-_R4-Pad1_ GND Net-_R5-Pad2_ APPS1 Net-_U1-Pad14_ MCP6004		
R1  Net-_R1-Pad1_ APPS1 1000		
R2  Net-_R2-Pad1_ APPS2 1000		
R4  Net-_R4-Pad1_ Net-_R1-Pad1_ 1000		
R3  GND Net-_R2-Pad1_ 1000		
U5  Net-_U5-Pad1_ Net-_R6-Pad2_ APPS1 +10V Net-_R8-Pad2_ APPS2 Net-_U5-Pad7_ Net-_U5-Pad8_ Net-_R10-Pad1_ APPS2 RTN_+5V_ MCP6004		
R11  +5V Net-_R11-Pad2_ 4750		
R13  Net-_R12-Pad2_ GND 4750		
R12  Net-_R11-Pad2_ Net-_R12-Pad2_ 500		
U6  Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U5-Pad1_ Net-_U5-Pad7_ Net-_U5-Pad8_ ? VSS Net-_U1-Pad14_ ? ? ? ? ? VDD 4073		
U4  +24V GND +5V LM78M05CT		
U3  +24V GND RTN_+5V_ LM78M05CT		
U2  +24V GND +10V LM7810CT		
C1  APPS1 GND 0.1u		
C2  APPS2 GND 0.1u		
Q1  ? ? ? MMBF170		

.end
